library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.common_defs.all;

--! Processor control store

--! The control store is a ROM used to store the processor microprogram.
entity control_store is
  port (
    --! Address of the desired word
    address : in  ctrl_str_addr_type;
    --! Content of the addressed word
    word    : out ctrl_str_word_type
    );
end entity control_store;

--! Dataflow architecture for the control store
architecture dataflow of control_store is

  -- Constants
  constant words : ctrl_str_type := (
--BEGIN_WORDS_ENTRY0 => "000000110000000000000000000000001001",


0 => "000001001000000000000000000000001001",
1 => "010111100000000000000000000000001001",
2 => "000000000000000000000000000000000000",
3 => "000000000000000000000000000000000000",
4 => "000000000000000000000000000000000000",
5 => "000000000000000000000000000000000000",
6 => "000000111000001101010000001000000001",
7 => "000001000000001101010000001000010001",
8 => "000001001000000000000000000000001001",
9 => "000000000100001101010000001000010001",
10 => "000000000000000000000000000000000000",
11 => "000000000000000000000000000000000000",
12 => "000000000000000000000000000000000000",
13 => "000000000000000000000000000000000000",
14 => "000000000000000000000000000000000000",
15 => "000000000000000000000000000000000000",
16 => "000010001000001101010000010010000100",
17 => "000010010000001101010000001000010001",
18 => "000001001000000101000010000101000010",
19 => "000000000000000000000000000000000000",
20 => "000000000000000000000000000000000000",
21 => "000010110000000101001000000000000101",
22 => "000010111000001111000000000010100011",
23 => "000011000000001101010000010010000100",
24 => "000011001000001101010000001001010001",
25 => "000001001000000101000010000000000000",
26 => "000000000000000000000000000000000000",
27 => "000000000000000000000000000000000000",
28 => "000000000000000000000000000000000000",
29 => "000000000000000000000000000000000000",
30 => "000000000000000000000000000000000000",
31 => "000000000000000000000000000000000000",
32 => "000100001000001101010000001000010001",
33 => "000100010000100101001000000000000011",
34 => "000100011000000111001000000000000011",
35 => "000010111000001111000000000010100110",
36 => "000000000000000000000000000000000000",
37 => "000000000000000000000000000000000000",
38 => "000000000000000000000000000000000000",
39 => "000000000000000000000000000000000000",
40 => "000000000000000000000000000000000000",
41 => "000000000000000000000000000000000000",
42 => "000000000000000000000000000000000000",
43 => "000000000000000000000000000000000000",
44 => "000000000000000000000000000000000000",
45 => "000000000000000000000000000000000000",
46 => "000000000000000000000000000000000000",
47 => "000000000000000000000000000000000000",
48 => "000000000000000000000000000000000000",
49 => "000000000000000000000000000000000000",
50 => "000000000000000000000000000000000000",
51 => "000000000000000000000000000000000000",
52 => "000000000000000000000000000000000000",
53 => "000000000000000000000000000000000000",
54 => "000110111000000101001000000000000101",
55 => "000111000000001111000000000010000011",
56 => "000111001000000101000000000101000111",
57 => "000111010000001101100000010010100100",
58 => "000111011000001101010000001000010001",
59 => "000001001000000101000010000000000000",
60 => "000000000000000000000000000000000000",
61 => "000000000000000000000000000000000000",
62 => "000000000000000000000000000000000000",
63 => "000000000000000000000000000000000000",
64 => "000000000000000000000000000000000000",
65 => "000000000000000000000000000000000000",
66 => "000000000000000000000000000000000000",
67 => "000000000000000000000000000000000000",
68 => "000000000000000000000000000000000000",
69 => "000000000000000000000000000000000000",
70 => "000000000000000000000000000000000000",
71 => "000000000000000000000000000000000000",
72 => "000000000000000000000000000000000000",
73 => "000000000000000000000000000000000000",
74 => "000000000000000000000000000000000000",
75 => "000000000000000000000000000000000000",
76 => "000000000000000000000000000000000000",
77 => "000000000000000000000000000000000000",
78 => "000000000000000000000000000000000000",
79 => "000000000000000000000000000000000000",
80 => "000000000000000000000000000000000000",
81 => "000000000000000000000000000000000000",
82 => "000000000000000000000000000000000000",
83 => "000000000000000000000000000000000000",
84 => "000000000000000000000000000000000000",
85 => "000000000000000000000000000000000000",
86 => "000000000000000000000000000000000000",
87 => "001011000000001101010000010010000100",
88 => "000001001000000101000000000101000111",
89 => "001011010000001101100000010010100100",
90 => "001011011000000000000000000000001001",
91 => "000001001000000101000010000000000000",
92 => "001011101000001101100000000010100100",
93 => "001011110000001101010000010010000100",
94 => "001011111000000101001000000000000111",
95 => "000001001000001111110010000101000000",
96 => "000000000000000000000000000000000000",
97 => "000000000000000000000000000000000000",
98 => "000000000000000000000000000000000000",
99 => "000000000000000000000000000000000000",
100 => "000000000000000000000000000000000000",
101 => "001100110000001101100000010010100100",
102 => "001100111000000101001000000000000111",
103 => "000001001000001111000010000101000000",
104 => "000000000000000000000000000000000000",
105 => "000000000000000000000000000000000000",
106 => "000000000000000000000000000000000000",
107 => "000000000000000000000000000000000000",
108 => "000000000000000000000000000000000000",
109 => "000000000000000000000000000000000000",
110 => "000000000000000000000000000000000000",
111 => "000000000000000000000000000000000000",
112 => "000000000000000000000000000000000000",
113 => "000000000000000000000000000000000000",
114 => "000000000000000000000000000000000000",
115 => "000000000000000000000000000000000000",
116 => "000000000000000000000000000000000000",
117 => "000000000000000000000000000000000000",
118 => "000000000000000000000000000000000000",
119 => "000000000000000000000000000000000000",
120 => "000000000000000000000000000000000000",
121 => "000000000000000000000000000000000000",
122 => "000000000000000000000000000000000000",
123 => "000000000000000000000000000000000000",
124 => "000000000000000000000000000000000000",
125 => "000000000000000000000000000000000000",
126 => "001111111000001101100000010010100100",
127 => "010000000000000101001000000000000111",
128 => "000001001000000011000010000101000000",
129 => "000000000000000000000000000000000000",
130 => "000000000000000000000000000000000000",
131 => "000000000000000000000000000000000000",
132 => "010000101000000101001000000000000101",
133 => "010000110000001111000000000010100011",
134 => "010000111000001101010000001000010001",
135 => "010001000000000101001000000000000000",
136 => "010001001000001101010000001000010001",
137 => "000001001000001111000000000101000010",
138 => "000000000000000000000000000000000000",
139 => "000000000000000000000000000000000000",
140 => "000000000000000000000000000000000000",
141 => "000000000000000000000000000000000000",
142 => "000000000000000000000000000000000000",
143 => "000000000000000000000000000000000000",
144 => "000000000000000000000000000000000000",
145 => "000000000000000000000000000000000000",
146 => "000000000000000000000000000000000000",
147 => "000000000000000000000000000000000000",
148 => "000000000000000000000000000000000000",
149 => "000000000000000000000000000000000000",
150 => "000000000000000000000000000000000000",
151 => "000000000000000000000000000000000000",
152 => "000000000000000000000000000000000000",
153 => "010011010000001101100000010010100100",
154 => "010011011000000101000100000000000111",
155 => "010011100000000101000010000000000000",
156 => "000000110001000101000000000000001000",
157 => "010011110000001101100000010010100100",
158 => "010011111000000101000100000000000111",
159 => "010100000000000101000010000000000000",
160 => "000000110010000101000000000000001000",
161 => "010100010000001101100000010010100100",
162 => "010100011000001101100000010010000100",
163 => "010100100000000101001000000000100000",
164 => "010100101000000101000100000000000111",
165 => "010100110000000101000010000000000000",
166 => "000000110001001111110000000000001000",
167 => "010101000000001101100100000000000001",
168 => "010101001000001101010000001000010001",
169 => "010101010000100101001000000000000010",
170 => "010101011000000111001000000000000011",
171 => "010101100000001111000000001000011000",
172 => "000001001000000000000000000000001001",
173 => "010101110000000101000000010010100101",
174 => "010101111000000000000000000000001001",
175 => "010110000000000101000000100010100000",
176 => "010110001000001101010000000010000101",
177 => "010110010000000101000000001000110000",
178 => "010110011000000101000000000010000100",
179 => "010110100000000101000000100000000000",
180 => "010110101000000101000000000101000111",
181 => "000001001001001101100000000000000001",
182 => "010110111000001101100000010010100100",
183 => "010111000000000101001000000000000111",
184 => "000001001000000111000010000101000000",
185 => "010111010000001101010000001000010001",
186 => "010111011000100101001000000000000011",
187 => "010111100000000111001000000000000011",
188 => "010111101000001111000000000010100110",
189 => "010111110000001101010100000000000001",
190 => "010111111000000101000000001000010000",
191 => "011000000000001101010000001000010001",
192 => "011000001000100101001000000000000011",
193 => "011000010000000111001000000000000011",
194 => "011000011000001101010000001000010001",
195 => "011000100000001111110010000000000100",
196 => "011000101000001101010010000010000111",
197 => "011000110000001101010000001000010001",
198 => "011000111000100101001000000000000011",
199 => "011001000000000111001000000000000011",
200 => "011001001000001111010000000101000100",
201 => "011001010000000101000000010010000000",
202 => "011001011000000101000000000101001000",
203 => "011001100000001101010000010010000100",
204 => "011001101000000101000000000101000101",
205 => "011001110000001101010000001000010001",
206 => "000001001000000101000000100000000111",
207 => "100000000100001101010000001000010001",
208 => "000000000000000000000000000000000000",
209 => "000000000000000000000000000000000000",
210 => "000000000000000000000000000000000000",
211 => "000000000000000000000000000000000000",
212 => "000000000000000000000000000000000000",
213 => "000000000000000000000000000000000000",
214 => "000000000000000000000000000000000000",
215 => "000000000000000000000000000000000000",
216 => "000000000000000000000000000000000000",
217 => "000000000000000000000000000000000000",
218 => "000000000000000000000000000000000000",
219 => "000000000000000000000000000000000000",
220 => "000000000000000000000000000000000000",
221 => "000000000000000000000000000000000000",
222 => "000000000000000000000000000000000000",
223 => "000000000000000000000000000000000000",
224 => "000000000000000000000000000000000000",
225 => "000000000000000000000000000000000000",
226 => "000000000000000000000000000000000000",
227 => "000000000000000000000000000000000000",
228 => "000000000000000000000000000000000000",
229 => "000000000000000000000000000000000000",
230 => "000000000000000000000000000000000000",
231 => "000000000000000000000000000000000000",
232 => "000000000000000000000000000000000000",
233 => "000000000000000000000000000000000000",
234 => "000000000000000000000000000000000000",
235 => "000000000000000000000000000000000000",
236 => "000000000000000000000000000000000000",
237 => "000000000000000000000000000000000000",
238 => "000000000000000000000000000000000000",
239 => "000000000000000000000000000000000000",
240 => "000000000000000000000000000000000000",
241 => "000000000000000000000000000000000000",
242 => "000000000000000000000000000000000000",
243 => "000000000000000000000000000000000000",
244 => "000000000000000000000000000000000000",
245 => "000000000000000000000000000000000000",
246 => "000000000000000000000000000000000000",
247 => "000000000000000000000000000000000000",
248 => "000000000000000000000000000000000000",
249 => "000000000000000000000000000000000000",
250 => "000000000000000000000000000000000000",
251 => "000000000000000000000000000000000000",
252 => "000000000000000000000000000000000000",
253 => "000000000000000000000000000000000000",
254 => "000000000000000000000000000000000000",
255 => "000000000000000000000000000000000000",
256 => "000000000000000000000000000000000000",
257 => "000000000000000000000000000000000000",
258 => "000000000000000000000000000000000000",
259 => "000000000000000000000000000000000000",
260 => "000000000000000000000000000000000000",
261 => "000000000000000000000000000000000000",
262 => "010101000000001101100100000000010001",
263 => "000000000000000000000000000000000000",
264 => "000000000000000000000000000000000000",
265 => "100001001000000000000000000000001001",
266 => "000000000000000000000000000000000000",
267 => "000000000000000000000000000000000000",
268 => "000000000000000000000000000000000000",
269 => "000000000000000000000000000000000000",
270 => "000000000000000000000000000000000000",
271 => "000000000000000000000000000000000000",
272 => "000000000000000000000000000000000000",
273 => "000000000000000000000000000000000000",
274 => "000000000000000000000000000000000000",
275 => "000000000000000000000000000000000000",
276 => "000000000000000000000000000000000000",
277 => "100010110000001101010000001000010001",
278 => "100010111000100101001000000000000011",
279 => "100011000000000111001000000000000011",
280 => "000010111000001111000000000010100101",
281 => "000000000000000000000000000000000000",
282 => "000000000000000000000000000000000000",
283 => "000000000000000000000000000000000000",
284 => "000000000000000000000000000000000000",
285 => "000000000000000000000000000000000000",
286 => "000000000000000000000000000000000000",
287 => "000000000000000000000000000000000000",
288 => "000000000000000000000000000000000000",
289 => "000000000000000000000000000000000000",
290 => "000000000000000000000000000000000000",
291 => "000000000000000000000000000000000000",
292 => "000000000000000000000000000000000000",
293 => "000000000000000000000000000000000000",
294 => "000000000000000000000000000000000000",
295 => "000000000000000000000000000000000000",
296 => "000000000000000000000000000000000000",
297 => "000000000000000000000000000000000000",
298 => "000000000000000000000000000000000000",
299 => "000000000000000000000000000000000000",
300 => "000000000000000000000000000000000000",
301 => "000000000000000000000000000000000000",
302 => "000000000000000000000000000000000000",
303 => "000000000000000000000000000000000000",
304 => "000000000000000000000000000000000000",
305 => "000000000000000000000000000000000000",
306 => "000000000000000000000000000000000000",
307 => "000000000000000000000000000000000000",
308 => "000000000000000000000000000000000000",
309 => "000000000000000000000000000000000000",
310 => "100110111000001101010000001000010001",
311 => "100111000000100101001000000000000011",
312 => "100111001000000111001000000000000011",
313 => "000111000000001111000000000010000101",
314 => "000000000000000000000000000000000000",
315 => "000000000000000000000000000000000000",
316 => "000000000000000000000000000000000000",
317 => "000000000000000000000000000000000000",
318 => "000000000000000000000000000000000000",
319 => "000000000000000000000000000000000000",
320 => "000000000000000000000000000000000000",
321 => "000000000000000000000000000000000000",
322 => "000000000000000000000000000000000000",
323 => "000000000000000000000000000000000000",
324 => "000000000000000000000000000000000000",
325 => "000000000000000000000000000000000000",
326 => "000000000000000000000000000000000000",
327 => "000000000000000000000000000000000000",
328 => "000000000000000000000000000000000000",
329 => "000000000000000000000000000000000000",
330 => "000000000000000000000000000000000000",
331 => "000000000000000000000000000000000000",
332 => "000000000000000000000000000000000000",
333 => "000000000000000000000000000000000000",
334 => "000000000000000000000000000000000000",
335 => "000000000000000000000000000000000000",
336 => "000000000000000000000000000000000000",
337 => "000000000000000000000000000000000000",
338 => "000000000000000000000000000000000000",
339 => "000000000000000000000000000000000000",
340 => "000000000000000000000000000000000000",
341 => "000000000000000000000000000000000000",
342 => "000000000000000000000000000000000000",
343 => "000000000000000000000000000000000000",
344 => "000000000000000000000000000000000000",
345 => "000000000000000000000000000000000000",
346 => "000000000000000000000000000000000000",
347 => "000000000000000000000000000000000000",
348 => "000000000000000000000000000000000000",
349 => "000000000000000000000000000000000000",
350 => "000000000000000000000000000000000000",
351 => "000000000000000000000000000000000000",
352 => "000000000000000000000000000000000000",
353 => "000000000000000000000000000000000000",
354 => "000000000000000000000000000000000000",
355 => "000000000000000000000000000000000000",
356 => "000000000000000000000000000000000000",
357 => "000000000000000000000000000000000000",
358 => "000000000000000000000000000000000000",
359 => "000000000000000000000000000000000000",
360 => "000000000000000000000000000000000000",
361 => "000000000000000000000000000000000000",
362 => "000000000000000000000000000000000000",
363 => "000000000000000000000000000000000000",
364 => "000000000000000000000000000000000000",
365 => "000000000000000000000000000000000000",
366 => "000000000000000000000000000000000000",
367 => "000000000000000000000000000000000000",
368 => "000000000000000000000000000000000000",
369 => "000000000000000000000000000000000000",
370 => "000000000000000000000000000000000000",
371 => "000000000000000000000000000000000000",
372 => "000000000000000000000000000000000000",
373 => "000000000000000000000000000000000000",
374 => "000000000000000000000000000000000000",
375 => "000000000000000000000000000000000000",
376 => "000000000000000000000000000000000000",
377 => "000000000000000000000000000000000000",
378 => "000000000000000000000000000000000000",
379 => "000000000000000000000000000000000000",
380 => "000000000000000000000000000000000000",
381 => "000000000000000000000000000000000000",
382 => "000000000000000000000000000000000000",
383 => "000000000000000000000000000000000000",
384 => "000000000000000000000000000000000000",
385 => "000000000000000000000000000000000000",
386 => "000000000000000000000000000000000000",
387 => "000000000000000000000000000000000000",
388 => "000000000000000000000000000000000000",
389 => "000000000000000000000000000000000000",
390 => "000000000000000000000000000000000000",
391 => "000000000000000000000000000000000000",
392 => "000000000000000000000000000000000000",
393 => "000000000000000000000000000000000000",
394 => "000000000000000000000000000000000000",
395 => "000000000000000000000000000000000000",
396 => "000000000000000000000000000000000000",
397 => "000000000000000000000000000000000000",
398 => "000000000000000000000000000000000000",
399 => "000000000000000000000000000000000000",
400 => "000000000000000000000000000000000000",
401 => "000000000000000000000000000000000000",
402 => "000000000000000000000000000000000000",
403 => "000000000000000000000000000000000000",
404 => "000000000000000000000000000000000000",
405 => "000000000000000000000000000000000000",
406 => "000000000000000000000000000000000000",
407 => "000000000000000000000000000000000000",
408 => "000000000000000000000000000000000000",
409 => "000000000000000000000000000000000000",
410 => "000000000000000000000000000000000000",
411 => "000000000000000000000000000000000000",
412 => "000000000000000000000000000000000000",
413 => "000000000000000000000000000000000000",
414 => "000000000000000000000000000000000000",
415 => "000000000000000000000000000000000000",
416 => "000000000000000000000000000000000000",
417 => "000000000000000000000000000000000000",
418 => "000000000000000000000000000000000000",
419 => "000000000000000000000000000000000000",
420 => "000000000000000000000000000000000000",
421 => "000000000000000000000000000000000000",
422 => "000000000000000000000000000000000000",
423 => "000000000000000000000000000000000000",
424 => "000000000000000000000000000000000000",
425 => "000000000000000000000000000000000000",
426 => "000000000000000000000000000000000000",
427 => "000000000000000000000000000000000000",
428 => "000000000000000000000000000000000000",
429 => "000000000000000000000000000000000000",
430 => "000000000000000000000000000000000000",
431 => "000000000000000000000000000000000000",
432 => "000000000000000000000000000000000000",
433 => "000000000000000000000000000000000000",
434 => "000000000000000000000000000000000000",
435 => "000000000000000000000000000000000000",
436 => "000000000000000000000000000000000000",
437 => "000000000000000000000000000000000000",
438 => "000000000000000000000000000000000000",
439 => "000000000000000000000000000000000000",
440 => "000000000000000000000000000000000000",
441 => "000000000000000000000000000000000000",
442 => "000000000000000000000000000000000000",
443 => "000000000000000000000000000000000000",
444 => "000000000000000000000000000000000000",
445 => "000000000000000000000000000000000000",
446 => "000000000000000000000000000000000000",
447 => "000000000000000000000000000000000000",
448 => "000000000000000000000000000000000000",
449 => "000000000000000000000000000000000000",
450 => "000000000000000000000000000000000000",
451 => "000000000000000000000000000000000000",
452 => "000000000000000000000000000000000000",
453 => "000000000000000000000000000000000000",
454 => "000000000000000000000000000000000000",
455 => "000000000000000000000000000000000000",
456 => "000000000000000000000000000000000000",
457 => "000000000000000000000000000000000000",
458 => "000000000000000000000000000000000000",
459 => "000000000000000000000000000000000000",
460 => "000000000000000000000000000000000000",
461 => "000000000000000000000000000000000000",
462 => "000000000000000000000000000000000000",
463 => "000000000000000000000000000000000000",
464 => "000000000000000000000000000000000000",
465 => "000000000000000000000000000000000000",
466 => "000000000000000000000000000000000000",
467 => "000000000000000000000000000000000000",
468 => "000000000000000000000000000000000000",
469 => "000000000000000000000000000000000000",
470 => "000000000000000000000000000000000000",
471 => "000000000000000000000000000000000000",
472 => "000000000000000000000000000000000000",
473 => "000000000000000000000000000000000000",
474 => "000000000000000000000000000000000000",
475 => "000000000000000000000000000000000000",
476 => "000000000000000000000000000000000000",
477 => "000000000000000000000000000000000000",
478 => "000000000000000000000000000000000000",
479 => "000000000000000000000000000000000000",
480 => "000000000000000000000000000000000000",
481 => "000000000000000000000000000000000000",
482 => "000000000000000000000000000000000000",
483 => "000000000000000000000000000000000000",
484 => "000000000000000000000000000000000000",
485 => "000000000000000000000000000000000000",
486 => "000000000000000000000000000000000000",
487 => "000000000000000000000000000000000000",
488 => "000000000000000000000000000000000000",
489 => "000000000000000000000000000000000000",
490 => "000000000000000000000000000000000000",
491 => "000000000000000000000000000000000000",
492 => "000000000000000000000000000000000000",
493 => "000000000000000000000000000000000000",
494 => "000000000000000000000000000000000000",
495 => "000000000000000000000000000000000000",
496 => "000000000000000000000000000000000000",
497 => "000000000000000000000000000000000000",
498 => "000000000000000000000000000000000000",
499 => "000000000000000000000000000000000000",
500 => "000000000000000000000000000000000000",
501 => "000000000000000000000000000000000000",
502 => "000000000000000000000000000000000000",
503 => "000000000000000000000000000000000000",
504 => "000000000000000000000000000000000000",
505 => "000000000000000000000000000000000000",
506 => "000000000000000000000000000000000000",
507 => "000000000000000000000000000000000000",
508 => "000000000000000000000000000000000000",
509 => "000000000000000000000000000000000000",
510 => "000000000000000000000000000000000000",
511 => "000000000000000000000000000000000000",

others => (others => '0')
--END_WORDS_ENTRY
    );

begin  -- architecture dataflow

  word <= words(to_integer(unsigned(address)));

end architecture dataflow;